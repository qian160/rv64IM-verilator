// virtual address -> physical address
module mmu(
    input   [38:0]  sv39_va_i,

    output  [38:0]  sv39_va_o,
    output  [55:0]  sv39_pa_o


);

endmodule

module tlb();

endmodule