module div(
    // todo
);

endmodule